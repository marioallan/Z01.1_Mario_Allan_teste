module and_verilog(

	input a, b,
	output c
);
	
	and(c, a, b);

endmodule
