module dut(

 input vint,
 output vout
 );

assign vout = vint;
 
endmodule
